module tb_ball_absolute_top();

endmodule


module d220324_dat_main();
    initial begin
        $display("d220324_dat_main module s");
        #200;
        $finish();

    end
endmodule