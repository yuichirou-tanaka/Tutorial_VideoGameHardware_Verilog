module tb_TestModule();
    d220324_dat_main d220324_dat_main_0();

    initial begin
        $display("test module s");
    end
endmodule